module second;

initial begin
$display("hello1");
$display("hello2");
end

endmodule
